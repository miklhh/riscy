--
-- Riscy RISC-V arithmetic and logic unit
-- Author: Mikael Henriksson (2023)
--

library ieee, work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.riscy_conf.all;

entity riscy_alu is

end entity riscy_alu;
